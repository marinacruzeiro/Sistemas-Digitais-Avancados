LIBRARY	IEEE;
USE IEEE.std_logic_1164.all;

PACKAGE type_array2 IS

	TYPE array_reg IS ARRAY (31 DOWNTO 0) OF STD_LOGIC_VECTOR (7 DOWNTO 0);

END type_array2;